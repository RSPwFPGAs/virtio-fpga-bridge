`include "dma_transaction_for_queue_notify.v"
